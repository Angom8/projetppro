Niveau3:1,Niveau1:2,Niveau4:3,Niveau5:0,Niveau3:0,Test:0#
