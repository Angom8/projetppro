VOID:0#
