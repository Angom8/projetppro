Niveau3:0,Niveau1:0#
